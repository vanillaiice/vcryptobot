module config

fn test_config() {
	println(new())
}
